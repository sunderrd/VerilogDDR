/*
 * --GRAPHICS MODULE--
 * directs graphics from the note positions to the vga controller
 */

module graphics(clk, rst);





endmodule